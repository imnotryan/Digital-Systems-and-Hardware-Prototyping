`timescale 1ns / 1ps


module tb_test_Systolic_Array();
    
    reg clk;
    reg start; 
    reg reset;
    reg [7:0] a00, a01, a02, a10, a11, a12, a20, a21, a22; // each a00, a01, etc is a register that is 8 bits long 
    reg [7:0] b00, b01, b02, b10, b11, b12, b20, b21, b22; // each b00, b01, etc is a register that is 8 bits long
    
    wire done;
    wire [7:0] M1_out, M2_out, M3_out, M4_out, M5_out, M6_out, M7_out, M8_out, M9_out;
    
    always #5 clk = ~clk;
    
    test_Systolic_Matrix uut( clk, reset, start, 
                a00, a01, a02, a10, a11, a12, a20, a21, a22, 
                b00, b01, b02, b10, b11, b12, b20, b21, b22,
                //make sure the above wires/ports are identicaly
                
                //You can choose not to have below wires/ports in your design
                M1_out, M2_out, M3_out, M4_out, M5_out, M6_out, M7_out, M8_out, M9_out, 
                done);
initial begin
    //input inputs here!
clk = 0;
reset = 1;
	
	// TEST SET 1
//        a00 = 8'b00110000; a01 = 8'b00110000; a02 = 8'b00110000;    //  1    1    1
//        a10 = 8'b00110000; a11 = 8'b00110000; a12 = 8'b00110000;    //  1    1    1
//        a20 = 8'b00110000; a21 = 8'b00110000; a22 = 8'b00110000;    //  1    1    1
    
//        b00 = 8'b00110000; b01 = 8'b00110000; b02 = 8'b00110000;    //  1    1    1
//        b10 = 8'b00110000; b11 = 8'b00110000; b12 = 8'b00110000;    //  1    1    1
//        b20 = 8'b00110000; b21 = 8'b00110000; b22 = 8'b00110000;    //  1    1    1
        
////        c00 = 8'b01001000; c01 = 8'b01001000; c02 = 8'b01001000;    //  3     3     3
////        c10 = 8'b01001000; c11 = 8'b01001000; c12 = 8'b01001000;    //  3     3     3
////        c20 = 8'b01001000; c01 = 8'b01001000; c02 = 8'b01001000;    //  3     3     3

//        #10
//        reset = 0;
//        #100
//        start = 1;

//        #200
//        reset = 1;
//        start = 0;

	// TEST SET 2
//        a00 = 8'b00110000; a01 = 8'b00110000; a02 = 8'b00110000;    //  1    1    1
//        a10 = 8'b00110000; a11 = 8'b00110000; a12 = 8'b00110000;    //  1    1    1
//        a20 = 8'b00110000; a21 = 8'b00110000; a22 = 8'b00110000;    //  1    1    1
    
//        b00 = 8'b00110000; b01 = 8'b10100000; b02 = 8'b00110000;    //  1     -0.5      1
//        b10 = 8'b10111000; b11 = 8'b01000000; b12 = 8'b10111000;    //  -1.5    2     -1.5
//        b20 = 8'b00110000; b21 = 8'b10100000; b22 = 8'b00110000;    //  1     -0.5       1
        
////        c00 = 8'b00100000; c01 = 8'b00110000; c02 = 8'b00100000;    //  0.5     1     0.5
////        c10 = 8'b00100000; c11 = 8'b00110000; c12 = 8'b00100000;    //  0.5     1     0.5
////        c20 = 8'b00100000; c21 = 8'b00110000; c22 = 8'b00100000;    //  0.5     1     0.5    

//        #10
//        reset = 0;
//        #100
//        start = 1;

//        #200
//        reset = 1;
//        start = 0;

	// TEST SET 3
	  a00 = 8'b00000000; a01 = 8'b00110000; a02 = 8'b00110000;    //  0    1    1
        a10 = 8'b00110000; a11 = 8'b00000000; a12 = 8'b00110000;    //  1    0    1
        a20 = 8'b00110000; a21 = 8'b00110000; a22 = 8'b00000000;    //  1    1    0
    
        b00 = 8'b00110000; b01 = 8'b10100000; b02 = 8'b00110000;    //  1     -0.5      1
        b10 = 8'b10111000; b11 = 8'b01000000; b12 = 8'b10111000;    //  -1.5    2     -1.5
        b20 = 8'b00110000; b21 = 8'b10100000; b22 = 8'b00110000;    //  1     -0.5       1
        
//        c00 = 8'b10100000; c01 = 8'b00111000; c02 = 8'b10100000;    //  -0.5     1.5     -0.5
//        c10 = 8'b01000000; c11 = 8'b10110000; c12 = 8'b01000000;    //    2     -1       2
//        c20 = 8'b10100000; c01 = 8'b00111000; c02 = 8'b10100000;    //  -0.5     1.5     -0.5 

        #10
        reset = 0;
        #100
        start = 1;


     
end
endmodule
